* C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab3\Q2\q2.sch

* Schematics Version 8.0 - July 1997
* Fri May 14 11:13:49 2010



** Analysis setup **
.OP 
.LIB "C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab3\Q2\q2.lib"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "q2.net"
.INC "q2.als"


.probe


.END
