* C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab4\Q1\Q1.sch

* Schematics Version 8.0 - July 1997
* Fri Jul 02 13:57:10 2010



** Analysis setup **
.tran 20ns 10ms
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "Q1.net"
.INC "Q1.als"


.probe


.END
