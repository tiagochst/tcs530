* C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab4\Q2\Q2.sch

* Schematics Version 8.0 - July 1997
* Sat Jul 03 09:01:38 2010



** Analysis setup **
.DC LIN V_V3 -10 10 0.1 
.tran 20ns 10ms
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "Q2.net"
.INC "Q2.als"


.probe


.END
