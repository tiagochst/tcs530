* C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab3\Q2\q2a.sch

* Schematics Version 8.0 - July 1997
* Fri May 21 22:25:11 2010



** Analysis setup **
.ac DEC 10 100 100000k
.tran/OP 20ns 100ms SKIPBP
.OP 
.LIB "C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab3\Q2\q2.lib"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib "C:\Users\Tiago\Desktop\EE530\pspice\tcs530\Lab3\Q1\q1.lib"
.lib "nom.lib"

.INC "q2a.net"
.INC "q2a.als"


.probe


.END
